`ifndef SPECS_VH
`define SPECS_VH

// supported opcodes
`define OP_SUM  3'b000
`define OP_SUB  3'b001
`define OP_AND  3'b010
`define OP_XOR  3'b011
`define OP_NOP  3'b100

// supported cpu bit width
`define WORD 8

`endif // SPECS_VH